package Test;

interface Ifc_type;
  method Action collatz_submit(Int#(64) n);
  method ActionValue#(Int#(64)) collatz_get();
endinterface: Ifc_type

interface Ifc_type;
  method Action collatz_submit(Int#(64) n);
  method ActionValue#(Int#(64)) collatz_get();
endinterface: Ifc_type


endpackage: Test
